    entity SNM_BO is
        port (

            p in : bit;
            soma out : natural 
            fd
            
        );
    end entity SNM_BO;

    architecture design of SNM_BO is
        
    begin
        
        
        
    end architecture design;