    entity SNM_BO is
        port (

            state in : bit;
            sum out : natural 
            
            
        );
    end entity SNM_BO;

    architecture design of SNM_BO is
        
    begin
        
        
        
    end architecture design;