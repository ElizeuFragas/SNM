    entity SNM_BO is
        port (

        	type tipo_estado is (A, B, C, D, E);
            state in : tipo_estado;
            sum out : interger; 
            
            
        );
    end entity SNM_BO;

    architecture behave of SNM_BO is
        
    begin
        
        
        
    end architecture behave;