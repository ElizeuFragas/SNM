entity SNM_BC is
    port (

        p in : bit;
        
        
    );
end entity SNM_BC;