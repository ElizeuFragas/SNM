entity SNM is
    port (
        
    );
end entity SNM;

architecture design of SNM is
    
begin
    
    
    
end architecture design;